`timescale 1ns / 1ps

module port_match#PORT_NUM#_#MODULEID#(port_no,final_mv,test_clk);
parameter w=#COMPSIZE#;
parameter n=#NO_OF_RULES#;
input [w-1:0] port_no;
input test_clk;
output reg [n-1:0] final_mv;

